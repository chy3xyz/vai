// vai.agent.coordination - 高级协调模式
// 实现 Map-Reduce、投票共识、管道处理等协作模式
module agent

import time
import json
import skills
import protocol { new_event_message }

// MapReduceJob Map-Reduce 作业
pub struct MapReduceJob {
pub:
	id          string
	description string
	input_data  []map[string]skills.Value // 输入数据集
	mapper      ?fn (map [string]skills.Value) map[string]skills.Value  // 映射函数
	reducer     ?fn ([]map[string]skills.Value) map[string]skills.Value // 归约函数
	num_workers int = 3
}

// MapReduceResult Map-Reduce 结果
pub struct MapReduceResult {
pub:
	job_id         string
	mapped_results []map[string]skills.Value
	final_result   map[string]skills.Value
	took_ms        i64
}

// 执行 Map-Reduce 作业
pub fn (mut h AgentHub) execute_mapreduce(job MapReduceJob) !MapReduceResult {
	start := time.now()

	// 获取工作节点
	workers := h.get_agents_by_role(.worker)
	if workers.len == 0 {
		return error('no worker agents available')
	}

	// Map 阶段
	mut mapped_results := []map[string]skills.Value{}
	mut map_tasks := []Task{}

	for i, data in job.input_data {
		task := Task{
			id:          '${job.id}_map_${i}'
			type_:       'map'
			description: 'Map task ${i} for job ${job.id}'
			input_data:  {
				'data':   data
				'mapper': 'custom'
			}
			priority:    0
		}
		map_tasks << task
	}

	// 分发 Map 任务
	for i, task in map_tasks {
		worker_idx := i % workers.len
		_ := workers[worker_idx]

		// 提交任务到工作节点
		h.task_queue <- task

		// 等待结果（简化实现）
		// 实际应该异步收集结果
	}

	// 等待所有 Map 任务完成
	time.sleep(2 * time.second)

	// Reduce 阶段
	reduce_task := Task{
		id:          '${job.id}_reduce'
		type_:       'reduce'
		description: 'Reduce task for job ${job.id}'
		input_data:  {
			'mapped': skills.Value(mapped_results)
		}
		priority:    1
	}

	// 查找规划者或协调者执行 Reduce
	planners := h.get_agents_by_role(.planner)
	if planners.len > 0 {
		_ := planners[0]
		h.task_queue <- reduce_task
	}

	took := time.since(start)

	return MapReduceResult{
		job_id:         job.id
		mapped_results: mapped_results
		final_result:   map[string]skills.Value{}
		took_ms:        took.milliseconds()
	}
}

// VotingProposal 投票提案
pub struct VotingProposal {
pub:
	id          string
	topic       string
	options     []string
	timeout_sec int = 60
}

// Vote 投票
pub struct Vote {
pub:
	proposal_id string
	voter_id    string
	choice      string
	reason      string
	timestamp   time.Time
}

// VotingResult 投票结果
pub struct VotingResult {
pub:
	proposal_id string
	votes       map[string][]string // 选项 -> 投票者列表
	winner      string
	consensus   f32 // 共识度 0-1
}

// 发起投票
pub fn (mut h AgentHub) initiate_voting(proposal VotingProposal) !VotingResult {
	// 获取所有 Agent
	agents := h.list_agents()

	mut votes := map[string]Vote{}

	// 向每个 Agent 发送投票请求
	for ag_info in agents {
		vote_request := new_event_message('vote_request', {
			'proposal': json.encode(proposal)
		})

		h.route_message('hub', ag_info.id, vote_request)!
	}

	// 等待投票结果
	time.sleep(proposal.timeout_sec * time.second)

	// 统计结果
	mut vote_counts := map[string][]string{}
	for _, vote in votes {
		if vote.choice !in vote_counts {
			vote_counts[vote.choice] = []
		}
		vote_counts[vote.choice] << vote.voter_id
	}

	// 找出获胜选项
	mut winner := ''
	mut max_votes := 0
	for option, voters in vote_counts {
		if voters.len > max_votes {
			max_votes = voters.len
			winner = option
		}
	}

	// 计算共识度
	consensus := if agents.len > 0 { f32(max_votes) / f32(agents.len) } else { 0.0 }

	return VotingResult{
		proposal_id: proposal.id
		votes:       vote_counts
		winner:      winner
		consensus:   consensus
	}
}

// PipelineStage 管道阶段
pub struct PipelineStage {
pub:
	id          string
	name        string
	processor   string // Agent ID
	input_type  string
	output_type string
}

// Pipeline 处理管道
pub struct Pipeline {
pub:
	id     string
	name   string
	stages []PipelineStage
	hub    &AgentHub
}

// 创建管道
pub fn (mut h AgentHub) create_pipeline(name string, stages []PipelineStage) !Pipeline {
	// 验证所有处理器都存在
	for stage in stages {
		if stage.processor !in h.agents {
			return error('processor not found: ${stage.processor}')
		}
	}

	return Pipeline{
		id:     generate_task_id()
		name:   name
		stages: stages
		hub:    &h
	}
}

// 执行管道处理
pub fn (mut p Pipeline) process(data map[string]skills.Value) !map[string]skills.Value {
	mut current_data := data.clone()

	for stage in p.stages {
		// 创建处理任务
		task := Task{
			id:          '${p.id}_${stage.id}'
			type_:       'pipeline_stage'
			description: 'Pipeline stage: ${stage.name}'
			input_data:  current_data
			assigned_to: stage.processor
		}

		// 提交任务
		p.hub.task_queue <- task

		// 等待结果（简化实现）
		time.sleep(500 * time.millisecond)

		// 获取结果
		if res := p.hub.results[task.id] {
			if res.success {
				current_data = res.output.clone()
			} else {
				return error('pipeline stage ${stage.name} failed: ${res.error_msg}')
			}
		}
	}

	return current_data
}

// ConsensusBuilder 共识构建器
// 用于多 Agent 达成共识决策
pub struct ConsensusBuilder {
pub mut:
	hub          &AgentHub
	participants []string
	rounds       int = 3
}

// 创建共识构建器
pub fn new_consensus_builder(hub &AgentHub, participants []string) ConsensusBuilder {
	return ConsensusBuilder{
		hub:          hub
		participants: participants
		rounds:       3
	}
}

// 执行共识流程
pub fn (mut cb ConsensusBuilder) reach_consensus(topic string, initial_proposal string) !string {
	mut current_proposal := initial_proposal

	for round := 0; round < cb.rounds; round++ {
		// TODO: collect feedbacks from participants

		// 收集反馈
		for participant_id in cb.participants {
			feedback_task := Task{
				id:          'consensus_${round}_${participant_id}'
				type_:       'feedback'
				description: 'Provide feedback on: ${current_proposal}'
				input_data:  {
					'proposal': skills.Value(current_proposal)
					'topic':    skills.Value(topic)
					'round':    skills.Value(i64(round))
				}
				assigned_to: participant_id
			}

			cb.hub.task_queue <- feedback_task
		}

		// 等待反馈
		time.sleep(2 * time.second)

		// 整合反馈生成新提案
		// 简化：直接返回当前提案
		if round == cb.rounds - 1 {
			return current_proposal
		}
	}

	return current_proposal
}

// LoadBalancer 负载均衡器
pub struct LoadBalancer {
pub mut:
	hub      &AgentHub
	strategy LoadBalanceStrategy = .least_connections
}

// 负载均衡策略
pub enum LoadBalanceStrategy {
	round_robin
	least_connections
	weighted_response_time
	capability_based
}

// 选择 Agent
pub fn (mut lb LoadBalancer) select_agent(task Task) ?&BaseAgent {
	match lb.strategy {
		.round_robin {
			workers := lb.hub.get_agents_by_role(.worker)
			if workers.len > 0 {
				idx := time.now().second % workers.len
				return workers[idx]
			}
		}
		.least_connections {
			mut min_load := 999999
			mut selected := ?&BaseAgent(none)

			for _, ag_info in lb.hub.agents {
				// 简化：使用状态作为负载指标
				load := if ag_info.agent_status == .busy { 1 } else { 0 }
				if load < min_load {
					min_load = load
					selected = unsafe { ag_info }
				}
			}
			return selected
		}
		.capability_based {
			// 选择能力最匹配的 Agent
			mut best_score := -1
			mut selected := ?&BaseAgent(none)

			for _, mut ag_info in lb.hub.agents {
				score := lb.calculate_capability_score(mut ag_info, task)
				if score > best_score {
					best_score = score
					selected = unsafe { ag_info }
				}
			}
			return selected
		}
		else {}
	}

	return none
}

// 计算能力匹配分数
fn (mut lb LoadBalancer) calculate_capability_score(mut ag BaseAgent, task Task) int {
	mut score := 0
	caps := ag.capabilities()
	_ := caps

	for req_cap in task.required_caps {
		if req_cap in caps {
			score += 10
		}
	}

	return score
}

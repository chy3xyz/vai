// vai.cli - 本地控制台/调试工具 (简化版)
module cli

import os
import term
import time

// CLI 命令行接口
@[heap]
pub struct CLI {
	pub mut:
		name           string
		version        string
		commands       map[string]Command
		prompt         string = 'vai> '
		history_file   string
		running        bool
}

// Command 命令接口
pub interface Command {
	name() string
	description() string
	aliases() []string
	execute(args []string, mut ctx Context) !
}

// Context 命令上下文
pub struct Context {
	pub mut:
		app_data map[string]voidptr
}

// BaseCommand 基础命令实现
pub struct BaseCommand {
	pub:
		cmd_name        string
		cmd_description string
		cmd_aliases     []string
}

pub fn (c BaseCommand) name() string {
	return c.cmd_name
}

pub fn (c BaseCommand) description() string {
	return c.cmd_description
}

pub fn (c BaseCommand) aliases() []string {
	return c.cmd_aliases
}

// 创建 CLI
pub fn new_cli(name string, version string) &CLI {
	return &CLI{
		name: name
		version: version
		commands: map[string]Command{}
		history_file: os.join_path(os.home_dir(), '.${name}_history')
	}
}

// 注册命令
pub fn (mut c CLI) register(cmd Command) {
	c.commands[cmd.name()] = cmd
	for alias in cmd.aliases() {
		c.commands[alias] = cmd
	}
}

// 运行 CLI
pub fn (mut c CLI) run() {
	c.running = true
	c.print_banner()

	for c.running {
		print(c.prompt)
		input := os.input('')
		line := input.trim_space()

		if line.len == 0 {
			continue
		}

		c.execute(line) or {
			println(term.red('Error: ${err}'))
		}
	}
}

// 执行命令
pub fn (mut c CLI) execute(line string) ! {
	parts := line.split(' ')
	if parts.len == 0 {
		return
	}

	cmd_name := parts[0]
	args := if parts.len > 1 { parts[1..] } else { []string{} }

	if cmd := c.commands[cmd_name] {
		mut ctx := Context{
			app_data: map[string]voidptr{}
		}
		cmd.execute(args, mut ctx)!
	} else {
		return error('unknown command: ${cmd_name}. Type "help" for available commands.')
	}
}

// 停止 CLI
pub fn (c &CLI) stop() {
	// 使用 unsafe 块来修改 running 状态
	// 这是因为 Command 接口要求 execute 方法使用不可变接收器
	unsafe {
		mut mutable_c := c
		mutable_c.running = false
	}
}

// 打印 Banner
fn (c &CLI) print_banner() {
	println('')
	println(term.cyan('╔════════════════════════════════════════╗'))
	println(term.cyan('║') + '  ${term.bold(c.name)} v${c.version}${' '.repeat(35 - c.name.len - c.version.len)}' + term.cyan('║'))
	println(term.cyan('║') + '  V AI Infrastructure Console${' '.repeat(22)}' + term.cyan('║'))
	println(term.cyan('╚════════════════════════════════════════╝'))
	println('')
	println('Type "help" for available commands, "quit" to exit.')
	println('')
}

// HelpCommand 帮助命令
pub struct HelpCommand {
	BaseCommand
	pub mut:
		cli_ptr &CLI
}

pub fn new_help_command(cli_ptr &CLI) HelpCommand {
	return HelpCommand{
		BaseCommand: BaseCommand{
			cmd_name: 'help'
			cmd_description: 'Show help information'
			cmd_aliases: ['h', '?']
		}
		cli_ptr: cli_ptr
	}
}

pub fn (c HelpCommand) execute(args []string, mut ctx Context) ! {
	if args.len > 0 {
		cmd_name := args[0]
		if cmd := c.cli_ptr.commands[cmd_name] {
			println('')
			println(term.bold('Command: ') + cmd.name())
			println(term.bold('Description: ') + cmd.description())
			aliases := cmd.aliases()
			if aliases.len > 0 {
				println(term.bold('Aliases: ') + aliases.join(', '))
			}
			println('')
		} else {
			return error('unknown command: ${cmd_name}')
		}
	} else {
		println('')
		println(term.bold('Available commands:'))
		println('')

		mut unique_commands := map[string]Command{}
		for _, cmd in c.cli_ptr.commands {
			unique_commands[cmd.name()] = cmd
		}

		for _, cmd in unique_commands {
			name := term.green(cmd.name())
			padding := ' '.repeat(15 - cmd.name().len)
			println('  ${name}${padding}${cmd.description()}')
		}

		println('')
	}
}

// QuitCommand 退出命令
pub struct QuitCommand {
	BaseCommand
	pub mut:
		cli_ptr &CLI
}

pub fn new_quit_command(cli_ptr &CLI) QuitCommand {
	return QuitCommand{
		BaseCommand: BaseCommand{
			cmd_name: 'quit'
			cmd_description: 'Exit the CLI'
			cmd_aliases: ['exit', 'q']
		}
		cli_ptr: cli_ptr
	}
}

pub fn (c QuitCommand) execute(args []string, mut ctx Context) ! {
	println('Goodbye!')
	c.cli_ptr.stop()
}

// VersionCommand 版本命令
pub struct VersionCommand {
	BaseCommand
	pub mut:
		cli_ptr &CLI
}

pub fn new_version_command(cli_ptr &CLI) VersionCommand {
	return VersionCommand{
		BaseCommand: BaseCommand{
			cmd_name: 'version'
			cmd_description: 'Show version information'
			cmd_aliases: ['v']
		}
		cli_ptr: cli_ptr
	}
}

pub fn (c VersionCommand) execute(args []string, mut ctx Context) ! {
	println('${c.cli_ptr.name} v${c.cli_ptr.version}')
}

// StatusInfo 状态信息
pub struct StatusInfo {
	pub:
		uptime           time.Duration
		active_agents  int
		messages_processed int
		memory_usage   string
}

// StatusCommand 状态命令
pub struct StatusCommand {
	BaseCommand
	pub mut:
		get_status fn () StatusInfo = unsafe { nil }
}

pub fn new_status_command(get_status fn () StatusInfo) StatusCommand {
	return StatusCommand{
		BaseCommand: BaseCommand{
			cmd_name: 'status'
			cmd_description: 'Show system status'
			cmd_aliases: ['st']
		}
		get_status: get_status
	}
}

pub fn (c StatusCommand) execute(args []string, mut ctx Context) ! {
	status := c.get_status()

	println('')
	println(term.bold('System Status'))
	println('  Uptime:         ${status.uptime}')
	println('  Active Agents:  ${status.active_agents}')
	println('  Messages:       ${status.messages_processed}')
	println('  Memory Usage:   ${status.memory_usage}')
	println('')
}

// ClearCommand 清屏命令
pub struct ClearCommand {
	BaseCommand
}

pub fn new_clear_command() ClearCommand {
	return ClearCommand{
		BaseCommand: BaseCommand{
			cmd_name: 'clear'
			cmd_description: 'Clear the screen'
			cmd_aliases: ['cls']
		}
	}
}

pub fn (c ClearCommand) execute(args []string, mut ctx Context) ! {
	print('\x1b[2J\x1b[H')
}

// EchoCommand 回显命令（用于测试）
pub struct EchoCommand {
	BaseCommand
}

pub fn new_echo_command() EchoCommand {
	return EchoCommand{
		BaseCommand: BaseCommand{
			cmd_name: 'echo'
			cmd_description: 'Echo the input'
			cmd_aliases: []
		}
	}
}

pub fn (c EchoCommand) execute(args []string, mut ctx Context) ! {
	println(args.join(' '))
}

// OnboardCommand 初始化命令
pub struct OnboardCommand {
	BaseCommand
}

pub fn new_onboard_command() OnboardCommand {
	return OnboardCommand{
		BaseCommand: BaseCommand{
			cmd_name: 'onboard'
			cmd_description: 'Initialize VAI configuration and workspace'
			cmd_aliases: ['init', 'setup']
		}
	}
}

pub fn (c OnboardCommand) execute(args []string, mut ctx Context) ! {
	println('Initializing VAI...')
	
	// 这里会调用配置和工作区初始化
	// 实际实现会在集成阶段完成
	println('VAI initialized successfully!')
	println('Configuration: ~/.vai/config.json')
	println('Workspace: ~/.vai/workspace/')
}

// CronListCommand Cron 任务列表命令
pub struct CronListCommand {
	BaseCommand
	pub mut:
		get_cron_service fn () voidptr = unsafe { nil }
}

pub fn new_cron_list_command(get_cron_service fn () voidptr) CronListCommand {
	return CronListCommand{
		BaseCommand: BaseCommand{
			cmd_name: 'cron'
			cmd_description: 'List cron jobs'
			cmd_aliases: ['cron-list']
		}
		get_cron_service: get_cron_service
	}
}

pub fn (c CronListCommand) execute(args []string, mut ctx Context) ! {
	if args.len > 0 && args[0] == 'list' {
		println('Cron jobs:')
		// 实际实现会在集成阶段完成
		println('  (No cron jobs configured)')
	} else {
		println('Usage: cron list')
	}
}

// 注册默认命令
pub fn register_default_commands(mut c CLI, get_status fn () StatusInfo) {
	c.register(new_help_command(&c))
	c.register(new_quit_command(&c))
	c.register(new_version_command(&c))
	c.register(new_status_command(get_status))
	c.register(new_clear_command())
	c.register(new_echo_command())
	c.register(new_onboard_command())
}
